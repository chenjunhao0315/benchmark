// Benchmark "int2float_91" written by ABC on Thu Dec 19 15:11:37 2024

module int2float_91 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10,
    po0, po1, po2, po3, po4, po5, po6  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10;
  output po0, po1, po2, po3, po4, po5, po6;
  wire new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25,
    new_n26, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34,
    new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42,
    new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50,
    new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n58, new_n59,
    new_n60, new_n61, new_n62, new_n64, new_n65, new_n66, new_n67, new_n68,
    new_n69, new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76,
    new_n77, new_n78, new_n79, new_n80, new_n81, new_n82, new_n83, new_n84,
    new_n85, new_n86, new_n87, new_n88, new_n89, new_n90, new_n91, new_n92,
    new_n93, new_n94, new_n96, new_n97, new_n98, new_n99, new_n100,
    new_n101, new_n103, new_n104, new_n105, new_n106, new_n107;
  assign new_n19 = ~pi07 & ~pi08;
  assign new_n20 = ~pi09 & ~pi10;
  assign new_n21 = new_n19 & new_n20;
  assign new_n22 = pi03 & new_n21;
  assign new_n23 = pi02 & pi06;
  assign new_n24 = new_n22 & new_n23;
  assign new_n25 = pi04 & pi05;
  assign new_n26 = new_n24 & new_n25;
  assign po6 = ~new_n21 | new_n26;
  assign new_n28 = ~pi06 & ~po6;
  assign new_n29 = ~pi01 & new_n28;
  assign new_n30 = ~pi07 & ~new_n22;
  assign new_n31 = pi10 & new_n30;
  assign new_n32 = pi06 & ~po6;
  assign new_n33 = ~pi10 & ~new_n32;
  assign new_n34 = pi05 & ~po6;
  assign new_n35 = ~pi09 & ~new_n34;
  assign new_n36 = new_n33 & new_n35;
  assign new_n37 = ~pi04 & new_n36;
  assign new_n38 = ~new_n31 & ~new_n37;
  assign new_n39 = ~new_n29 & new_n38;
  assign new_n40 = pi02 & ~po6;
  assign new_n41 = ~pi06 & ~new_n40;
  assign new_n42 = ~pi08 & ~new_n28;
  assign new_n43 = new_n36 & new_n42;
  assign new_n44 = ~pi03 & new_n43;
  assign new_n45 = pi00 & new_n28;
  assign new_n46 = pi05 & new_n33;
  assign new_n47 = ~new_n45 & ~new_n46;
  assign new_n48 = ~new_n44 & ~new_n47;
  assign new_n49 = new_n39 & new_n48;
  assign new_n50 = ~new_n41 & new_n49;
  assign new_n51 = ~new_n36 & ~new_n50;
  assign new_n52 = ~new_n30 & new_n50;
  assign new_n53 = ~pi04 & ~po6;
  assign new_n54 = ~new_n52 & ~new_n53;
  assign new_n55 = new_n36 & ~new_n54;
  assign new_n56 = ~pi03 & ~new_n23;
  assign po3 = ~new_n55 | ~new_n56;
  assign new_n58 = ~new_n42 & ~new_n53;
  assign new_n59 = new_n52 & new_n58;
  assign new_n60 = po3 & new_n59;
  assign new_n61 = ~new_n36 & new_n60;
  assign new_n62 = ~new_n52 & ~new_n58;
  assign po5 = ~new_n36 | new_n60;
  assign new_n64 = ~new_n24 & ~po5;
  assign new_n65 = ~new_n62 & new_n64;
  assign new_n66 = new_n30 & new_n65;
  assign new_n67 = ~new_n61 & ~new_n66;
  assign new_n68 = new_n33 & new_n67;
  assign new_n69 = new_n51 & new_n68;
  assign new_n70 = ~new_n41 & ~new_n52;
  assign new_n71 = new_n51 & new_n70;
  assign new_n72 = ~new_n43 & ~new_n71;
  assign new_n73 = new_n47 & new_n72;
  assign new_n74 = ~new_n44 & ~new_n73;
  assign new_n75 = new_n39 & new_n74;
  assign new_n76 = ~new_n69 & ~new_n75;
  assign new_n77 = new_n39 & new_n76;
  assign new_n78 = new_n74 & new_n76;
  assign new_n79 = new_n29 & new_n55;
  assign new_n80 = new_n41 & new_n65;
  assign new_n81 = ~new_n24 & new_n42;
  assign new_n82 = new_n47 & new_n81;
  assign new_n83 = ~new_n80 & ~new_n82;
  assign new_n84 = ~new_n79 & new_n83;
  assign new_n85 = new_n35 & new_n84;
  assign new_n86 = ~new_n62 & ~new_n85;
  assign new_n87 = new_n67 & new_n86;
  assign new_n88 = ~new_n22 & ~new_n40;
  assign new_n89 = ~new_n87 & new_n88;
  assign new_n90 = ~new_n24 & ~new_n72;
  assign new_n91 = ~new_n89 & new_n90;
  assign new_n92 = new_n69 & new_n75;
  assign new_n93 = ~new_n91 & ~new_n92;
  assign new_n94 = ~new_n78 & new_n93;
  assign po0 = new_n77 | ~new_n94;
  assign new_n96 = new_n54 & ~new_n76;
  assign new_n97 = ~new_n84 & ~new_n96;
  assign new_n98 = new_n85 & new_n96;
  assign new_n99 = new_n30 & new_n69;
  assign new_n100 = ~new_n52 & ~new_n99;
  assign new_n101 = ~new_n98 & new_n100;
  assign po1 = ~new_n97 & new_n101;
  assign new_n103 = new_n36 & new_n70;
  assign new_n104 = ~new_n66 & new_n103;
  assign new_n105 = ~new_n33 & ~new_n35;
  assign new_n106 = ~new_n87 & ~new_n105;
  assign new_n107 = ~new_n104 & new_n106;
  assign po2 = new_n98 | ~new_n107;
  assign po4 = new_n65 | ~new_n68;
endmodule


